module practica_11 ( 
	a,
	b,
	s_r,
	s_i,
	l_b,
	s
	) ;

input [2:0] a;
input [2:0] b;
input  s_r;
input  s_i;
inout  l_b;
inout [2:0] s;
