module sumador_restador ( 
	a,
	b,
	s_r,
	s_i,
	c_o,
	s
	) ;

input [2:0] a;
input [2:0] b;
input  s_r;
input  s_i;
inout  c_o;
inout [2:0] s;
