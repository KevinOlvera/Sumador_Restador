module bcd_3_bits ( 
	i,
	o
	) ;

input [4:0] i;
inout [9:0] o;
