module practica_11 ( 
	a,
	b,
	ci,
	s_r,
	l_b,
	s
	) ;

input [3:0] a;
input [3:0] b;
input  ci;
input  s_r;
inout  l_b;
inout [3:0] s;
